module test;
  initial $display("Working!");
endmodule